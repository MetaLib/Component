* Simple LED Model
.subckt simpleLED 1 2
Dledx 1 2  DLed_test
.model Dled_test D (IS=8.6990E-18 RS=22.257 N=3.1999)
.ends